localparam    [2:0] addalu = 3'b000;
localparam    [2:0] subalu = 3'b001;
localparam    [2:0] andalu = 3'b010;